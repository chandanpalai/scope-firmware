--------------------------------------------------------------------------------
-- Engineer:       Ali Lown
--
-- Create Date:    19:38:54 08/14/2011
-- Module Name:    inputBoard - Behavioral
-- Project Name:   USB Digital Oscilloscope
-- Target Devices: xc3s50a(n)
-- Description:    Handles communications to/from the input boards uC's.
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity simplefifo is
  Port ( DATAIN : in STD_LOGIC_VECTOR(15 downto 0);
         WRCLK : in STD_LOGIC;
         DATAOUT : out STD_LOGIC_VECTOR(15 downto 0);
         RDCLK : in STD_LOGIC;
         FULL : out STD_LOGIC;
         EMPTY : out STD_LOGIC;
         RESET : in STD_LOGIC
       );
end simplefifo;

architecture Behavioral of simplefifo is

  constant maxcount : integer := 4;
  signal wrcount, rdcount : integer range 0 to maxcount := 0;
  type data_type is array((maxcount-1) downto 0) of std_logic_vector(15 downto 0);
  signal data : data_type;
  signal full_out, empty_out : std_logic;
begin
  FLAGS: process (RESET, wrcount, rdcount)
  begin
    if RESET = '1' then
      empty_out <= '1';
      full_out <= '0';
    end if;

    if wrcount > 0 then
      empty_out <= '0';
    else
      empty_out <= '1';
    end if;

    if wrcount = (maxcount-1) then
      full_out <= '1';
    else
      full_out <= '0';
    end if;
  end process;

  EMPTY <= empty_out;
  FULL <= full_out;

  WRITE: process (RESET, DATAIN, WRCLK, wrcount, full_out)
  begin
    if RESET = '1' then
      wrcount <= 0;
    else
      if WRCLK'event and WRCLK = '1' then
        if full_out = '0' then
          data(wrcount) <= DATAIN;
          wrcount <= wrcount + 1;
        end if;
      end if;
    end if;
  end process;

  READ: process (RESET, RDCLK, rdcount, empty_out)
  begin
    if RESET = '1' then
      rdcount <= 0;
    else
      if RDCLK'event and RDCLK = '1' then
        if empty_out = '0' then
          DATAOUT <= data(rdcount);
          rdcount <= rdcount + 1;
          if rdcount = (maxcount-1) then
            rdcount <= 0;
          end if;
        end if;
      end if;
    end if;
  end process;
end Behavioral;
